`ifndef _SRAM_SVH_
`define _SRAM_SVH_


// These will be used to determine which
parameter SRAM_ADDR_WIDTH = 4;
parameter SRAM_DATA_WIDTH = 8;






